module core_top (
    input clk,    // Clock
    input rst_n,  // Asynchronous reset active low


    input
    output  [INSTR_ADDR_WIDTH-1 : 0] o_instr_addr,    // 取指地址

);

endmodule